`ifndef SLAVE_DRIVER_SV
`define SLAVE_DRIVER_SV

class slave_driver extends uvm_driver #(slave_item);

  `uvm_component_utils(slave_driver)

  virtual slave_if vif;
  
  // Slave Req and Slave Res objects
  slave_item req;
  slave_item res;

  extern function new(string name, uvm_component parent);
  extern function void build_phase(uvm_phase phase);

  // Methods run_phase and do_drive generated by setting driver_inc in file slave.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_drive();

endclass : slave_driver 


function slave_driver::new(string name, uvm_component parent);
  super.new(name, parent);
endfunction : new


function void slave_driver::build_phase(uvm_phase phase);
  if (!uvm_config_db #(virtual slave_if)::get(this, "" , "slave_vif", vif))
    `uvm_fatal(get_type_name(), "Could not get virtual slave_if");
endfunction : build_phase


task slave_driver::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)
  
  forever begin
   
   // Monitor Ready Signal
   seq_item_port.get_next_item(req);
   seq_item_port.item_done();
      
   	wait(vif.ready);
   		repeat(10) begin
   			seq_item_port.get_next_item(res);
   			seq_item_port.item_done();
   	
   			// Driver Sequence to DUT
   			@(posedge vif.clk);
   			vif.valid	<= res.valid;
   			vif.data	<= res.data;
      		end
      		
      		@(posedge vif.clk);
   		vif.valid	<= 0;
   		vif.data	<= 0;
   end
endtask : run_phase



`endif // SLAVE_DRIVER_SV

